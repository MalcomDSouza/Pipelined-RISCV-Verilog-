module adder(
input signed [31:0]a,
input signed [31:0]b,
output [31:0]out);


assign out = a+b;


endmodule